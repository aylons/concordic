aylons@aylons-yoga2.26349:1399051022